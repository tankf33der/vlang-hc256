module hc256
